--o controller gia xeirismo diakopwn, den exw
--tin paramikri idea pws tha ylopoiithei gia tin wra
